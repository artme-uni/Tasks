`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.03.2019 19:58:08
// Design Name: 
// Module Name: tb_muxer16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_muxer16();

    logic [15:0] in;
    logic [0:0] q;
    logic [3:0] sel;
    
    muxer16 DUT(
    .in(in),
    .q(q),
    .sel(sel)
    );
    
initial begin
    sel = 4'b0000; in = 16'b0000000000000001; #10;
    sel = 4'b0000; in = 16'b1111111111111110; #10;

    sel = 4'b0001; in = 16'b0000000000000010; #10;
    sel = 4'b0001; in = 16'b1111111111111101; #10;
    
    sel = 4'b0010; in = 16'b0000000000000100; #10;
    sel = 4'b0010; in = 16'b1111111111111011; #10;
    
    sel = 4'b0011; in = 16'b0000000000001000; #10;   
    sel = 4'b0011; in = 16'b1111111111110111; #10;    
    
    sel = 4'b0100; in = 16'b0000000000010000; #10;      
    sel = 4'b0100; in = 16'b1111111111101111; #10;  
    
    sel = 4'b0101; in = 16'b0000000000100000; #10;
    sel = 4'b0101; in = 16'b1111111111011111; #10;
    
    sel = 4'b0110; in = 16'b0000000001000000; #10;
    sel = 4'b0110; in = 16'b1111111110111111; #10;
    
    sel = 4'b0111; in = 16'b0000000010000000; #10;
    sel = 4'b0111; in = 16'b1111111101111111; #10;
    
    sel = 4'b1000; in = 16'b0000000100000000; #10;
    sel = 4'b1000; in = 16'b1111111011111111; #10;
    
    sel = 4'b1001; in = 16'b0000001000000000; #10;
    sel = 4'b1001; in = 16'b1111110111111111; #10;
    
    sel = 4'b1010; in = 16'b0000010000000000; #10;
    sel = 4'b1010; in = 16'b1111101111111111; #10;
    
    sel = 4'b1011; in = 16'b0000100000000000; #10;
    sel = 4'b1011; in = 16'b1111011111111111; #10;
    
    sel = 4'b1100; in = 16'b0001000000000000; #10;
    sel = 4'b1100; in = 16'b1110111111111111; #10;
    
    sel = 4'b1101; in = 16'b0010000000000000; #10;
    sel = 4'b1101; in = 16'b1101111111111111; #10;
    
    sel = 4'b1110; in = 16'b0100000000000000; #10;
    sel = 4'b1110; in = 16'b1011111111111111; #10;
    
    sel = 4'b1111; in = 16'b1000000000000000; #10;
    sel = 4'b1111; in = 16'b0111111111111111; #10;
    
    $finish;
    end;
    
endmodule
