`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.03.2019 11:15:10
// Design Name: 
// Module Name: tb_sum
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_sum();

    logic [63:0] a;
    logic [63:0] b;
    logic cin;
    logic cout;
    logic [63:0] s;

sum64 DUT(.a(a), .b(b), .cin(cin), .s(s), .cout(cout));

initial begin
    {cin, a, b} = 129'b001010101010101010101010101010101010101010101010101010101010101011010101010101010101010101010101010101010101010101010101010101010; #10;
    {cin, a, b} = 129'b010101010101010101010101010101010101010101010101010101010101010100101010101010101010101010101010101010101010101010101010101010101; #10;
    
    {cin, a, b} = 129'b001010101010101010101010101010101010101010101010101010101010101011010101010101010101010101010101010101010101010101010101010101010; #10;
    {cin, a, b} = 129'b010101010101010101010101010101010101010101010101010101010101010100101010101010101010101010101010101010101010101010101010101010101; #10;    

    end
    
$finish;
end;

endmodule

